library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE CONVWERTER IS

	FUNCTION INT_TO_ASCI (A:INTEGER) RETURN STD_LOGIC_VECTOR;
	PROCEDURE SPLIT_NUMBER (SIGNAL NUMBER: IN INTEGER; SIGNAL DIGIT1,DIGIT2,DIGIT3: OUT INTEGER RANGE 0 TO 9);

END CONVWERTER;

PACKAGE BODY CONVWERTER IS

	FUNCTION INT_TO_ASCI (A:INTEGER) RETURN STD_LOGIC_VECTOR IS
	VARIABLE RESULT: STD_LOGIC_VECTOR(7 downto 0);
	BEGIN

	CASE A IS 
		WHEN 0 => RESULT:="00110000";
		WHEN 1 => RESULT:="00110001";
		WHEN 2 => RESULT:="00110010";
		WHEN 3 => RESULT:="00110011";
		WHEN 4 => RESULT:="00110100";
		WHEN 5 => RESULT:="00110101";
		WHEN 6 => RESULT:="00110110";
		WHEN 7 => RESULT:="00110111";
		WHEN 8 => RESULT:="00111000";
		WHEN 9 => RESULT:="00111001";
		WHEN OTHERS => RESULT:=(OTHERS=>'0');
	END CASE;	
	RETURN RESULT;
	END INT_TO_ASCI;
----------------------------------------------------------------------------------------------

	PROCEDURE SPLIT_NUMBER (SIGNAL NUMBER: IN INTEGER; SIGNAL DIGIT1,DIGIT2,DIGIT3: OUT INTEGER RANGE 0 TO 9) IS
		VARIABLE TEMP: INTEGER RANGE 0 TO 9999;
		VARIABLE D1: INTEGER RANGE 0 TO 9;
		VARIABLE D2: INTEGER RANGE 0 TO 9;
		VARIABLE D3: INTEGER RANGE 0 TO 9;
		BEGIN

		TEMP:=NUMBER;
		
		IF(TEMP>99)THEN
			D3:=TEMP/100;
			TEMP:=TEMP-D3*100;
		ELSE
			D3:=0;
		END IF;
		
		IF(TEMP>9)THEN
			D2:=TEMP/10;
			TEMP:=TEMP-D2*10;
		ELSE
			D2:=0;
		END IF;
		
		D1:=TEMP;

		DIGIT1<=D1;
		DIGIT2<=D2;
		DIGIT3<=D3;
	
	END SPLIT_NUMBER;
END CONVWERTER;